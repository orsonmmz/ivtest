// Copyright (c) 2015 CERN
// Maciej Suminski <maciej.suminski@cern.ch>
//
// This source code is free software; you can redistribute it
// and/or modify it in source code form under the terms of the GNU
// General Public License as published by the Free Software
// Foundation; either version 2 of the License, or (at your option)
// any later version.
//
// This program is distributed in the hope that it will be useful,
// but WITHOUT ANY WARRANTY; without even the implied warranty of
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
// GNU General Public License for more details.
//
// You should have received a copy of the GNU General Public License
// along with this program; if not, write to the Free Software
// Foundation, Inc., 59 Temple Place - Suite 330, Boston, MA 02111-1307, USA


// Test for time scaling functions $ivlh_time_from_def & $ivlh_time_to_def

module mod(input wire time a);
  timeunit 1us;
  timeprecision 1ps;

  always @(a) begin
    #($ivlh_time_from_def(a) + 1ns) $display("this message should appear first (time=%t)", $time());
  end
endmodule

module mod_test;
  timeunit 1ns;
  timeprecision 1fs;

  time a;
  mod dut(a);

  initial begin
    a <= $ivlh_time_to_def(3ns);
    #(5ns) $display("this message should appear second (time=%t)", $time());
  end
endmodule

